.title Basic Amplifier
.include '180nm_bulk.txt'
Vdd vdd 0 1.8V
R1 vdd out 50kOhm
M1 out in 0 0 nmos l=90nm w=1um
Vin in 0 DC 0.3V AC 1

.op
.end