.title Single-Stage Amplifier with PMOS Diode-Connected Load
Vdd Vdd 0 1.8
Vin in 0 DC 0.15 AC 1
M1 out in 0 0 nm l=90n w=1u
M2 out out Vdd Vdd pm l=90n w=1u
.model nm nmos level=14 version=4.8.1
.model pm nmos level=14 version=4.8.1
.op
.end