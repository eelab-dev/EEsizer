.title Basic circuit
.include '180nm_bulk.txt'
mp1 out a vdd vdd pmos L=90n W=10u   
mp2 out b vdd vdd pmos L=90n W=10u  
mn1 out a n1  0 nmos L=90n W=10u   
mn2 n1  b 0 0 nmos L=90n W=10u   

Vdd vdd 0 DC 1.8
Va a 0 pulse (0 1.8 0 0.1n 0.1n 25n 50n)
Vb b 0 pulse (0 1.8 0 0.1n 0.1n 40n 80n)

.end